module OpLUT
(
);

	parameter INSTRUCTION_CNT	10
	parameter OP_BITS		6
	parameter FUNC_BITS		6
	reg [INSTRUCTION_CNT:0] 	rom	[0:OP_BITS+FUNC_BITS];

	initial
		
	end

endmodule

1001_0000000000001010   //PC= 4  addi $t1,$0,10
101011_01000_00000_0000000000000000   //PC= 8  sw $0,0($t0)
101011_01000_01001_0000000000000100   //PC=12  sw $t1,4($t0)
100011_01000_01101_0000000000000100   //PC=16  lw $t5,4($t0)
000000_01101_01001_01111_00000_100000 //PC=20  add $t7,$t5,$t1       (hazard!)  
001000_00000_01010_0000000000001101   //PC=24  addi $t2,$0,13        (stall 1 cycle)
000000_01001_01001_01011_00000_011000 //PC=28  mul $t3,$t1,$t1
000010_00000000000000000000001011     //PC=32  j Jump            
001000_01001_01001_0000000000000001   //PC=36  addi $t1,$t1,1        (flush)
001000_01001_01001_0000000000000001   //PC=40  addi $t1,$t1,1        
000000_01010_01001_01010_00000_100010 //PC=44  Jump: sub $t2,$t2,$t1
000000_01001_01010_01011_00000_100100 //PC=48  and $t3,$t1,$t2
000000_01010_01011_01100_00000_100101 //PC=52  or $t4,$t2,$t3

