module GeneralControl
(
);

endmodule
