module L1_Cache
(
);

endmodule
