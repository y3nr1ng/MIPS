module GeneralControl
(
	
);

endmodule
