module L1_Cache_Controller
(
);

endmodule
