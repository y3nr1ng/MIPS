module ForwardingUnit(
	input	[]	IDEX_Rs,
	input	[]	IDEX_Rt,
	input	[]	EXMEM_Rd,
	input	[]	MEMWB_Rd,
	output	[0:1]	ALUdata1_sel,
	output	[0:1]	ALUdata2_sel
);


endmodule