`include "LookupTable.v"

module ALUControl (
);

endmodule
